`timescale 1ns / 1ps

module mux16_test;

	// Inputs
	reg [15:0] X;
	reg [3:0] C;

	// Outputs
	wire Y;

	// Instantiate the Unit Under Test (UUT)
	mux16 uut (
		.X(X), 
		.C(C), 
		.Y(Y)
	);

	initial begin
		// X = 1110110010000011
		X = 16'b1110110010000011;
		C = 4'b0000;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b0001;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b0010;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b0011;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b0100;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b0101;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b0110;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b0111;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b1000;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b1001;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b1010;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b1011;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b1100;
		#100;
        
		X = 16'b1110110010000011;
		C = 4'b1101;
		#100;

		X = 16'b1110110010000011;
		C = 4'b1110;
		#100;
		
		X = 16'b1110110010000011;
		C = 4'b1111;
		#100;
		
		// X = 1001001110110001
		X = 16'b1001001110110001;
		C = 4'b0000;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b0001;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b0010;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b0011;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b0100;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b0101;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b0110;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b0111;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b1000;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b1001;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b1010;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b1011;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b1100;
		#100;
        
		X = 16'b1001001110110001;
		C = 4'b1101;
		#100;

		X = 16'b1001001110110001;
		C = 4'b1110;
		#100;
		
		X = 16'b1001001110110001;
		C = 4'b1111;
		#100;
	end
      
endmodule

